* Simulation of pv cell
*
.tran 0.01ms 5ms uic
.include pv.net

.control
set color0 = white
set color1 = black
run
plot i(vse) vs v(nv) v(nv)*i(vse)/40 vs v(nv)
.endc
